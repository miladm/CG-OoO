.param Nw=64
.param Nh=64
