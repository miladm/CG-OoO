** Parametrized NAND2

.subckt nand2 a b y vdd_l
mp1    y  a  vdd_l  vdd_l  pmos L=2 W='Wp'
mp2    y  b  vdd_l  vdd_l  pmos L=2 W='Wp'
mn1    y  a  n1     0      nmos L=2 W='Wn'
mn2    n1 b  0      0      nmos L=2 W='Wn'
.ends

** .subckt dut a y vdd_l
** x1     clk  inp  y      vdd_l  nand2
** .ends
