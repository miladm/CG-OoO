.param Wn=2398.87
.param Wp=7196.60
.param Wload=27508.178
.param Rload=55.776
.include "inv.ckt"
