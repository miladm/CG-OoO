.param Nw=166
.param Nh=64
