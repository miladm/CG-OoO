.param Nw=86
.param Nh=16
