.param Wn=22.72
.param Wp=68.15
.param Wload=170.797
.param Rload=2.688
.include "inv.ckt"
