.param Nw=66
.param Nh=4
