.param Wn=67.16
.param Wp=201.49
.param Wload=705.869
.param Rload=14.336
.include "inv.ckt"
