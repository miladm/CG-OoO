.param Wn3=6
.param Wn=2
.param Wp=2
