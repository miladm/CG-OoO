.param Wn=116.31
.param Wp=348.94
.param Wload=704.539
.param Rload=11.088
.include "inv.ckt"
