.param Wn=167.07
.param Wp=501.20
.param Wload=1836.071
.param Rload=28.896
.include "inv.ckt"
