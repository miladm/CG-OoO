.param Nw=32
.param Nh=4
